// Code your testbench here
// or browse Examples
module hello_world;
  initial begin
    $display("Hello, World! Welcome to my 60-Day Verilog Challenge!");
    $finish;
  end
endmodule

